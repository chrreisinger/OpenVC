a + b sll 1 <= c*d and not e 
