assert expr report "some string" severity ERROR;
