loop
  exit when expr1;
  next when expr2;
end loop;

