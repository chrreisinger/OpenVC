type rec is record
  a : integer;
  b : real;
end record;


