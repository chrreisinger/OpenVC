function sin (s : real) return real;
attribute foreign of sin [real return real] : function 
   is "java.lang.Math";
