variable a : myEnum;
a := myEnum'value("first");
report myEnum'image(a);


