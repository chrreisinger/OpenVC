if condition1 then
  target := expr1;
elsif condition2 then
  target := expr2;
... 
elsif conditionN
  target := exprN;
end if;
