with expression select
target := 
  expr1 when choiceList1,
  expr2 when choiceList2,
  ...
  exprN when choiceListN;
