if expr1 then
  statement1;
elsif expr2 then
  statement2;
else
  statement3;
end if;
