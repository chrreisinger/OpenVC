while expr loop 
     statement1; 
     statement2; 
end loop; 
