package body p is
  procedure proc(x : IntA) is 
  begin
  end;
  procedure proc(x : IntB) is 
  begin
  end;
end p;

