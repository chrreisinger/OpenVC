constant PI : real := 3.14159_26535_89793_23846;