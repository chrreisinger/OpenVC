target :=
  expr1 when condition1 else
  expr2 when condition2 else
  ... 
  exprN when conditionN;
