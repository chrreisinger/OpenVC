type myEnum is (first, second, third);

