case expression is
  when choiceList1 => target := expr1;
  when choiceList2 => target := expr2;
  ...
  when choiceListN => target := exprN;
end case;
