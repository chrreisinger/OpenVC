for i in 0 to 10 loop
  null;
end loop
