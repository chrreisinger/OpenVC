variable x : integer range 5 to 10;
x := expr; 


