for i in 10 downto 0 loop
  null;
end loop
